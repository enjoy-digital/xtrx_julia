-------------------------------------------------------------------------------
-- Title      : i2c waveform ROM for xtrx power init sequencer
-- Project    : 
-------------------------------------------------------------------------------
-- File       : xtrxinitrom.vhd
-- Author     : mazsi-on-xtrx <>
-- Company    : 
-- Created    : 2019-02-21
-- Last update: 2019-03-05
-- Platform   : 
-- Standard   : VHDL'93/02
-------------------------------------------------------------------------------
-- Description: generated by xtrxinitgen.py -- should map into a single BRAM
--
-- with extra registers on address input and data output
-------------------------------------------------------------------------------
-- Copyright (c) 2019 GPLv2 (no later versions)
-------------------------------------------------------------------------------
-- Revisions  :
-- Date        Author  Description
-- 2019-02-21  mazsi   Created
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;

entity xtrxinitrom is

  port (
    CLK : in  std_logic;
    A   : in  std_logic_vector(11 downto 0);
    Q   : out std_logic_vector(3 downto 0)  -- bus, scl, sda, check
    );

end entity xtrxinitrom;

architecture imp of xtrxinitrom is
  signal a1   : std_logic_vector(A'range);
  signal qpre : std_logic_vector(Q'range);
begin

  process (CLK)
  begin
    if CLK'event and CLK = '1' then

      a1 <= A;

      case a1 is
        -- reset bus 0: idle, start, stop, idle
        when x"000" => qpre <= "0110";
        when x"001" => qpre <= "0110";
        when x"002" => qpre <= "0110";
        when x"003" => qpre <= "0110";
        when x"004" => qpre <= "0110";
        when x"005" => qpre <= "0100";
        when x"006" => qpre <= "0100";
        when x"007" => qpre <= "0000";
        when x"008" => qpre <= "0000";
        when x"009" => qpre <= "0100";
        when x"00a" => qpre <= "0100";
        when x"00b" => qpre <= "0110";
        when x"00c" => qpre <= "0110";
        when x"00d" => qpre <= "0110";
        when x"00e" => qpre <= "0110";
        when x"00f" => qpre <= "0110";
        -- reset bus 1: idle, start, stop, idle
        when x"010" => qpre <= "1110";
        when x"011" => qpre <= "1110";
        when x"012" => qpre <= "1110";
        when x"013" => qpre <= "1110";
        when x"014" => qpre <= "1110";
        when x"015" => qpre <= "1100";
        when x"016" => qpre <= "1100";
        when x"017" => qpre <= "1000";
        when x"018" => qpre <= "1000";
        when x"019" => qpre <= "1100";
        when x"01a" => qpre <= "1100";
        when x"01b" => qpre <= "1110";
        when x"01c" => qpre <= "1110";
        when x"01d" => qpre <= "1110";
        when x"01e" => qpre <= "1110";
        when x"01f" => qpre <= "1110";
        -- PMICL: check OTP ID
        when x"100" => qpre <= "0110";
        when x"101" => qpre <= "0110";
        when x"102" => qpre <= "0110";
        when x"103" => qpre <= "0110";
        when x"104" => qpre <= "0110";
        when x"105" => qpre <= "0100";
        when x"106" => qpre <= "0100";
        when x"107" => qpre <= "0000";
        when x"108" => qpre <= "0010";
        when x"109" => qpre <= "0110";
        when x"10a" => qpre <= "0110";
        when x"10b" => qpre <= "0010";
        when x"10c" => qpre <= "0010";
        when x"10d" => qpre <= "0110";
        when x"10e" => qpre <= "0110";
        when x"10f" => qpre <= "0010";
        when x"110" => qpre <= "0000";
        when x"111" => qpre <= "0100";
        when x"112" => qpre <= "0100";
        when x"113" => qpre <= "0000";
        when x"114" => qpre <= "0000";
        when x"115" => qpre <= "0100";
        when x"116" => qpre <= "0100";
        when x"117" => qpre <= "0000";
        when x"118" => qpre <= "0000";
        when x"119" => qpre <= "0100";
        when x"11a" => qpre <= "0100";
        when x"11b" => qpre <= "0000";
        when x"11c" => qpre <= "0000";
        when x"11d" => qpre <= "0100";
        when x"11e" => qpre <= "0100";
        when x"11f" => qpre <= "0000";
        when x"120" => qpre <= "0000";
        when x"121" => qpre <= "0100";
        when x"122" => qpre <= "0100";
        when x"123" => qpre <= "0000";
        when x"124" => qpre <= "0000";
        when x"125" => qpre <= "0100";
        when x"126" => qpre <= "0100";
        when x"127" => qpre <= "0000";
        when x"128" => qpre <= "0001";
        when x"129" => qpre <= "0101";
        when x"12a" => qpre <= "0101";
        when x"12b" => qpre <= "0001";
        when x"12c" => qpre <= "0000";
        when x"12d" => qpre <= "0000";
        when x"12e" => qpre <= "0000";
        when x"12f" => qpre <= "0000";
        when x"130" => qpre <= "0000";
        when x"131" => qpre <= "0100";
        when x"132" => qpre <= "0100";
        when x"133" => qpre <= "0000";
        when x"134" => qpre <= "0000";
        when x"135" => qpre <= "0100";
        when x"136" => qpre <= "0100";
        when x"137" => qpre <= "0000";
        when x"138" => qpre <= "0000";
        when x"139" => qpre <= "0100";
        when x"13a" => qpre <= "0100";
        when x"13b" => qpre <= "0000";
        when x"13c" => qpre <= "0000";
        when x"13d" => qpre <= "0100";
        when x"13e" => qpre <= "0100";
        when x"13f" => qpre <= "0000";
        when x"140" => qpre <= "0000";
        when x"141" => qpre <= "0100";
        when x"142" => qpre <= "0100";
        when x"143" => qpre <= "0000";
        when x"144" => qpre <= "0000";
        when x"145" => qpre <= "0100";
        when x"146" => qpre <= "0100";
        when x"147" => qpre <= "0000";
        when x"148" => qpre <= "0000";
        when x"149" => qpre <= "0100";
        when x"14a" => qpre <= "0100";
        when x"14b" => qpre <= "0000";
        when x"14c" => qpre <= "0010";
        when x"14d" => qpre <= "0110";
        when x"14e" => qpre <= "0110";
        when x"14f" => qpre <= "0010";
        when x"150" => qpre <= "0001";
        when x"151" => qpre <= "0101";
        when x"152" => qpre <= "0101";
        when x"153" => qpre <= "0001";
        when x"154" => qpre <= "0010";
        when x"155" => qpre <= "0110";
        when x"156" => qpre <= "0100";
        when x"157" => qpre <= "0000";
        when x"158" => qpre <= "0010";
        when x"159" => qpre <= "0110";
        when x"15a" => qpre <= "0110";
        when x"15b" => qpre <= "0010";
        when x"15c" => qpre <= "0010";
        when x"15d" => qpre <= "0110";
        when x"15e" => qpre <= "0110";
        when x"15f" => qpre <= "0010";
        when x"160" => qpre <= "0000";
        when x"161" => qpre <= "0100";
        when x"162" => qpre <= "0100";
        when x"163" => qpre <= "0000";
        when x"164" => qpre <= "0000";
        when x"165" => qpre <= "0100";
        when x"166" => qpre <= "0100";
        when x"167" => qpre <= "0000";
        when x"168" => qpre <= "0000";
        when x"169" => qpre <= "0100";
        when x"16a" => qpre <= "0100";
        when x"16b" => qpre <= "0000";
        when x"16c" => qpre <= "0000";
        when x"16d" => qpre <= "0100";
        when x"16e" => qpre <= "0100";
        when x"16f" => qpre <= "0000";
        when x"170" => qpre <= "0000";
        when x"171" => qpre <= "0100";
        when x"172" => qpre <= "0100";
        when x"173" => qpre <= "0000";
        when x"174" => qpre <= "0010";
        when x"175" => qpre <= "0110";
        when x"176" => qpre <= "0110";
        when x"177" => qpre <= "0010";
        when x"178" => qpre <= "0001";
        when x"179" => qpre <= "0101";
        when x"17a" => qpre <= "0101";
        when x"17b" => qpre <= "0001";
        when x"17c" => qpre <= "0000";
        when x"17d" => qpre <= "0000";
        when x"17e" => qpre <= "0000";
        when x"17f" => qpre <= "0000";
        when x"180" => qpre <= "0011";
        when x"181" => qpre <= "0111";
        when x"182" => qpre <= "0111";
        when x"183" => qpre <= "0011";
        when x"184" => qpre <= "0011";
        when x"185" => qpre <= "0111";
        when x"186" => qpre <= "0111";
        when x"187" => qpre <= "0011";
        when x"188" => qpre <= "0011";
        when x"189" => qpre <= "0111";
        when x"18a" => qpre <= "0111";
        when x"18b" => qpre <= "0011";
        when x"18c" => qpre <= "0001";
        when x"18d" => qpre <= "0101";
        when x"18e" => qpre <= "0101";
        when x"18f" => qpre <= "0001";
        when x"190" => qpre <= "0001";
        when x"191" => qpre <= "0101";
        when x"192" => qpre <= "0101";
        when x"193" => qpre <= "0001";
        when x"194" => qpre <= "0001";
        when x"195" => qpre <= "0101";
        when x"196" => qpre <= "0101";
        when x"197" => qpre <= "0001";
        when x"198" => qpre <= "0001";
        when x"199" => qpre <= "0101";
        when x"19a" => qpre <= "0101";
        when x"19b" => qpre <= "0001";
        when x"19c" => qpre <= "0001";
        when x"19d" => qpre <= "0101";
        when x"19e" => qpre <= "0101";
        when x"19f" => qpre <= "0001";
        when x"1a0" => qpre <= "0010";
        when x"1a1" => qpre <= "0110";
        when x"1a2" => qpre <= "0110";
        when x"1a3" => qpre <= "0010";
        when x"1a4" => qpre <= "0000";
        when x"1a5" => qpre <= "0000";
        when x"1a6" => qpre <= "0000";
        when x"1a7" => qpre <= "0000";
        when x"1a8" => qpre <= "0000";
        when x"1a9" => qpre <= "0100";
        when x"1aa" => qpre <= "0100";
        when x"1ab" => qpre <= "0110";
        when x"1ac" => qpre <= "0110";
        when x"1ad" => qpre <= "0110";
        when x"1ae" => qpre <= "0110";
        when x"1af" => qpre <= "0110";
        -- PMICL: enable buck1
        when x"200" => qpre <= "0110";
        when x"201" => qpre <= "0110";
        when x"202" => qpre <= "0110";
        when x"203" => qpre <= "0110";
        when x"204" => qpre <= "0110";
        when x"205" => qpre <= "0100";
        when x"206" => qpre <= "0100";
        when x"207" => qpre <= "0000";
        when x"208" => qpre <= "0010";
        when x"209" => qpre <= "0110";
        when x"20a" => qpre <= "0110";
        when x"20b" => qpre <= "0010";
        when x"20c" => qpre <= "0010";
        when x"20d" => qpre <= "0110";
        when x"20e" => qpre <= "0110";
        when x"20f" => qpre <= "0010";
        when x"210" => qpre <= "0000";
        when x"211" => qpre <= "0100";
        when x"212" => qpre <= "0100";
        when x"213" => qpre <= "0000";
        when x"214" => qpre <= "0000";
        when x"215" => qpre <= "0100";
        when x"216" => qpre <= "0100";
        when x"217" => qpre <= "0000";
        when x"218" => qpre <= "0000";
        when x"219" => qpre <= "0100";
        when x"21a" => qpre <= "0100";
        when x"21b" => qpre <= "0000";
        when x"21c" => qpre <= "0000";
        when x"21d" => qpre <= "0100";
        when x"21e" => qpre <= "0100";
        when x"21f" => qpre <= "0000";
        when x"220" => qpre <= "0000";
        when x"221" => qpre <= "0100";
        when x"222" => qpre <= "0100";
        when x"223" => qpre <= "0000";
        when x"224" => qpre <= "0000";
        when x"225" => qpre <= "0100";
        when x"226" => qpre <= "0100";
        when x"227" => qpre <= "0000";
        when x"228" => qpre <= "0001";
        when x"229" => qpre <= "0101";
        when x"22a" => qpre <= "0101";
        when x"22b" => qpre <= "0001";
        when x"22c" => qpre <= "0000";
        when x"22d" => qpre <= "0000";
        when x"22e" => qpre <= "0000";
        when x"22f" => qpre <= "0000";
        when x"230" => qpre <= "0000";
        when x"231" => qpre <= "0100";
        when x"232" => qpre <= "0100";
        when x"233" => qpre <= "0000";
        when x"234" => qpre <= "0000";
        when x"235" => qpre <= "0100";
        when x"236" => qpre <= "0100";
        when x"237" => qpre <= "0000";
        when x"238" => qpre <= "0000";
        when x"239" => qpre <= "0100";
        when x"23a" => qpre <= "0100";
        when x"23b" => qpre <= "0000";
        when x"23c" => qpre <= "0000";
        when x"23d" => qpre <= "0100";
        when x"23e" => qpre <= "0100";
        when x"23f" => qpre <= "0000";
        when x"240" => qpre <= "0000";
        when x"241" => qpre <= "0100";
        when x"242" => qpre <= "0100";
        when x"243" => qpre <= "0000";
        when x"244" => qpre <= "0010";
        when x"245" => qpre <= "0110";
        when x"246" => qpre <= "0110";
        when x"247" => qpre <= "0010";
        when x"248" => qpre <= "0000";
        when x"249" => qpre <= "0100";
        when x"24a" => qpre <= "0100";
        when x"24b" => qpre <= "0000";
        when x"24c" => qpre <= "0000";
        when x"24d" => qpre <= "0100";
        when x"24e" => qpre <= "0100";
        when x"24f" => qpre <= "0000";
        when x"250" => qpre <= "0001";
        when x"251" => qpre <= "0101";
        when x"252" => qpre <= "0101";
        when x"253" => qpre <= "0001";
        when x"254" => qpre <= "0000";
        when x"255" => qpre <= "0000";
        when x"256" => qpre <= "0000";
        when x"257" => qpre <= "0000";
        when x"258" => qpre <= "0010";
        when x"259" => qpre <= "0110";
        when x"25a" => qpre <= "0110";
        when x"25b" => qpre <= "0010";
        when x"25c" => qpre <= "0000";
        when x"25d" => qpre <= "0100";
        when x"25e" => qpre <= "0100";
        when x"25f" => qpre <= "0000";
        when x"260" => qpre <= "0000";
        when x"261" => qpre <= "0100";
        when x"262" => qpre <= "0100";
        when x"263" => qpre <= "0000";
        when x"264" => qpre <= "0000";
        when x"265" => qpre <= "0100";
        when x"266" => qpre <= "0100";
        when x"267" => qpre <= "0000";
        when x"268" => qpre <= "0010";
        when x"269" => qpre <= "0110";
        when x"26a" => qpre <= "0110";
        when x"26b" => qpre <= "0010";
        when x"26c" => qpre <= "0000";
        when x"26d" => qpre <= "0100";
        when x"26e" => qpre <= "0100";
        when x"26f" => qpre <= "0000";
        when x"270" => qpre <= "0000";
        when x"271" => qpre <= "0100";
        when x"272" => qpre <= "0100";
        when x"273" => qpre <= "0000";
        when x"274" => qpre <= "0000";
        when x"275" => qpre <= "0100";
        when x"276" => qpre <= "0100";
        when x"277" => qpre <= "0000";
        when x"278" => qpre <= "0001";
        when x"279" => qpre <= "0101";
        when x"27a" => qpre <= "0101";
        when x"27b" => qpre <= "0001";
        when x"27c" => qpre <= "0000";
        when x"27d" => qpre <= "0000";
        when x"27e" => qpre <= "0000";
        when x"27f" => qpre <= "0000";
        when x"280" => qpre <= "0000";
        when x"281" => qpre <= "0100";
        when x"282" => qpre <= "0100";
        when x"283" => qpre <= "0110";
        when x"284" => qpre <= "0110";
        when x"285" => qpre <= "0110";
        when x"286" => qpre <= "0110";
        when x"287" => qpre <= "0110";
        -- PMICL: set buck1 to 3280 mV
        when x"300" => qpre <= "0110";
        when x"301" => qpre <= "0110";
        when x"302" => qpre <= "0110";
        when x"303" => qpre <= "0110";
        when x"304" => qpre <= "0110";
        when x"305" => qpre <= "0100";
        when x"306" => qpre <= "0100";
        when x"307" => qpre <= "0000";
        when x"308" => qpre <= "0010";
        when x"309" => qpre <= "0110";
        when x"30a" => qpre <= "0110";
        when x"30b" => qpre <= "0010";
        when x"30c" => qpre <= "0010";
        when x"30d" => qpre <= "0110";
        when x"30e" => qpre <= "0110";
        when x"30f" => qpre <= "0010";
        when x"310" => qpre <= "0000";
        when x"311" => qpre <= "0100";
        when x"312" => qpre <= "0100";
        when x"313" => qpre <= "0000";
        when x"314" => qpre <= "0000";
        when x"315" => qpre <= "0100";
        when x"316" => qpre <= "0100";
        when x"317" => qpre <= "0000";
        when x"318" => qpre <= "0000";
        when x"319" => qpre <= "0100";
        when x"31a" => qpre <= "0100";
        when x"31b" => qpre <= "0000";
        when x"31c" => qpre <= "0000";
        when x"31d" => qpre <= "0100";
        when x"31e" => qpre <= "0100";
        when x"31f" => qpre <= "0000";
        when x"320" => qpre <= "0000";
        when x"321" => qpre <= "0100";
        when x"322" => qpre <= "0100";
        when x"323" => qpre <= "0000";
        when x"324" => qpre <= "0000";
        when x"325" => qpre <= "0100";
        when x"326" => qpre <= "0100";
        when x"327" => qpre <= "0000";
        when x"328" => qpre <= "0001";
        when x"329" => qpre <= "0101";
        when x"32a" => qpre <= "0101";
        when x"32b" => qpre <= "0001";
        when x"32c" => qpre <= "0000";
        when x"32d" => qpre <= "0000";
        when x"32e" => qpre <= "0000";
        when x"32f" => qpre <= "0000";
        when x"330" => qpre <= "0000";
        when x"331" => qpre <= "0100";
        when x"332" => qpre <= "0100";
        when x"333" => qpre <= "0000";
        when x"334" => qpre <= "0000";
        when x"335" => qpre <= "0100";
        when x"336" => qpre <= "0100";
        when x"337" => qpre <= "0000";
        when x"338" => qpre <= "0000";
        when x"339" => qpre <= "0100";
        when x"33a" => qpre <= "0100";
        when x"33b" => qpre <= "0000";
        when x"33c" => qpre <= "0000";
        when x"33d" => qpre <= "0100";
        when x"33e" => qpre <= "0100";
        when x"33f" => qpre <= "0000";
        when x"340" => qpre <= "0010";
        when x"341" => qpre <= "0110";
        when x"342" => qpre <= "0110";
        when x"343" => qpre <= "0010";
        when x"344" => qpre <= "0010";
        when x"345" => qpre <= "0110";
        when x"346" => qpre <= "0110";
        when x"347" => qpre <= "0010";
        when x"348" => qpre <= "0000";
        when x"349" => qpre <= "0100";
        when x"34a" => qpre <= "0100";
        when x"34b" => qpre <= "0000";
        when x"34c" => qpre <= "0000";
        when x"34d" => qpre <= "0100";
        when x"34e" => qpre <= "0100";
        when x"34f" => qpre <= "0000";
        when x"350" => qpre <= "0001";
        when x"351" => qpre <= "0101";
        when x"352" => qpre <= "0101";
        when x"353" => qpre <= "0001";
        when x"354" => qpre <= "0000";
        when x"355" => qpre <= "0000";
        when x"356" => qpre <= "0000";
        when x"357" => qpre <= "0000";
        when x"358" => qpre <= "0010";
        when x"359" => qpre <= "0110";
        when x"35a" => qpre <= "0110";
        when x"35b" => qpre <= "0010";
        when x"35c" => qpre <= "0010";
        when x"35d" => qpre <= "0110";
        when x"35e" => qpre <= "0110";
        when x"35f" => qpre <= "0010";
        when x"360" => qpre <= "0010";
        when x"361" => qpre <= "0110";
        when x"362" => qpre <= "0110";
        when x"363" => qpre <= "0010";
        when x"364" => qpre <= "0010";
        when x"365" => qpre <= "0110";
        when x"366" => qpre <= "0110";
        when x"367" => qpre <= "0010";
        when x"368" => qpre <= "0010";
        when x"369" => qpre <= "0110";
        when x"36a" => qpre <= "0110";
        when x"36b" => qpre <= "0010";
        when x"36c" => qpre <= "0000";
        when x"36d" => qpre <= "0100";
        when x"36e" => qpre <= "0100";
        when x"36f" => qpre <= "0000";
        when x"370" => qpre <= "0010";
        when x"371" => qpre <= "0110";
        when x"372" => qpre <= "0110";
        when x"373" => qpre <= "0010";
        when x"374" => qpre <= "0010";
        when x"375" => qpre <= "0110";
        when x"376" => qpre <= "0110";
        when x"377" => qpre <= "0010";
        when x"378" => qpre <= "0001";
        when x"379" => qpre <= "0101";
        when x"37a" => qpre <= "0101";
        when x"37b" => qpre <= "0001";
        when x"37c" => qpre <= "0000";
        when x"37d" => qpre <= "0000";
        when x"37e" => qpre <= "0000";
        when x"37f" => qpre <= "0000";
        when x"380" => qpre <= "0000";
        when x"381" => qpre <= "0100";
        when x"382" => qpre <= "0100";
        when x"383" => qpre <= "0110";
        when x"384" => qpre <= "0110";
        when x"385" => qpre <= "0110";
        when x"386" => qpre <= "0110";
        when x"387" => qpre <= "0110";
        -- PMICL: disable buck0
        when x"400" => qpre <= "0110";
        when x"401" => qpre <= "0110";
        when x"402" => qpre <= "0110";
        when x"403" => qpre <= "0110";
        when x"404" => qpre <= "0110";
        when x"405" => qpre <= "0100";
        when x"406" => qpre <= "0100";
        when x"407" => qpre <= "0000";
        when x"408" => qpre <= "0010";
        when x"409" => qpre <= "0110";
        when x"40a" => qpre <= "0110";
        when x"40b" => qpre <= "0010";
        when x"40c" => qpre <= "0010";
        when x"40d" => qpre <= "0110";
        when x"40e" => qpre <= "0110";
        when x"40f" => qpre <= "0010";
        when x"410" => qpre <= "0000";
        when x"411" => qpre <= "0100";
        when x"412" => qpre <= "0100";
        when x"413" => qpre <= "0000";
        when x"414" => qpre <= "0000";
        when x"415" => qpre <= "0100";
        when x"416" => qpre <= "0100";
        when x"417" => qpre <= "0000";
        when x"418" => qpre <= "0000";
        when x"419" => qpre <= "0100";
        when x"41a" => qpre <= "0100";
        when x"41b" => qpre <= "0000";
        when x"41c" => qpre <= "0000";
        when x"41d" => qpre <= "0100";
        when x"41e" => qpre <= "0100";
        when x"41f" => qpre <= "0000";
        when x"420" => qpre <= "0000";
        when x"421" => qpre <= "0100";
        when x"422" => qpre <= "0100";
        when x"423" => qpre <= "0000";
        when x"424" => qpre <= "0000";
        when x"425" => qpre <= "0100";
        when x"426" => qpre <= "0100";
        when x"427" => qpre <= "0000";
        when x"428" => qpre <= "0001";
        when x"429" => qpre <= "0101";
        when x"42a" => qpre <= "0101";
        when x"42b" => qpre <= "0001";
        when x"42c" => qpre <= "0000";
        when x"42d" => qpre <= "0000";
        when x"42e" => qpre <= "0000";
        when x"42f" => qpre <= "0000";
        when x"430" => qpre <= "0000";
        when x"431" => qpre <= "0100";
        when x"432" => qpre <= "0100";
        when x"433" => qpre <= "0000";
        when x"434" => qpre <= "0000";
        when x"435" => qpre <= "0100";
        when x"436" => qpre <= "0100";
        when x"437" => qpre <= "0000";
        when x"438" => qpre <= "0000";
        when x"439" => qpre <= "0100";
        when x"43a" => qpre <= "0100";
        when x"43b" => qpre <= "0000";
        when x"43c" => qpre <= "0000";
        when x"43d" => qpre <= "0100";
        when x"43e" => qpre <= "0100";
        when x"43f" => qpre <= "0000";
        when x"440" => qpre <= "0000";
        when x"441" => qpre <= "0100";
        when x"442" => qpre <= "0100";
        when x"443" => qpre <= "0000";
        when x"444" => qpre <= "0000";
        when x"445" => qpre <= "0100";
        when x"446" => qpre <= "0100";
        when x"447" => qpre <= "0000";
        when x"448" => qpre <= "0010";
        when x"449" => qpre <= "0110";
        when x"44a" => qpre <= "0110";
        when x"44b" => qpre <= "0010";
        when x"44c" => qpre <= "0000";
        when x"44d" => qpre <= "0100";
        when x"44e" => qpre <= "0100";
        when x"44f" => qpre <= "0000";
        when x"450" => qpre <= "0001";
        when x"451" => qpre <= "0101";
        when x"452" => qpre <= "0101";
        when x"453" => qpre <= "0001";
        when x"454" => qpre <= "0000";
        when x"455" => qpre <= "0000";
        when x"456" => qpre <= "0000";
        when x"457" => qpre <= "0000";
        when x"458" => qpre <= "0010";
        when x"459" => qpre <= "0110";
        when x"45a" => qpre <= "0110";
        when x"45b" => qpre <= "0010";
        when x"45c" => qpre <= "0010";
        when x"45d" => qpre <= "0110";
        when x"45e" => qpre <= "0110";
        when x"45f" => qpre <= "0010";
        when x"460" => qpre <= "0000";
        when x"461" => qpre <= "0100";
        when x"462" => qpre <= "0100";
        when x"463" => qpre <= "0000";
        when x"464" => qpre <= "0000";
        when x"465" => qpre <= "0100";
        when x"466" => qpre <= "0100";
        when x"467" => qpre <= "0000";
        when x"468" => qpre <= "0010";
        when x"469" => qpre <= "0110";
        when x"46a" => qpre <= "0110";
        when x"46b" => qpre <= "0010";
        when x"46c" => qpre <= "0000";
        when x"46d" => qpre <= "0100";
        when x"46e" => qpre <= "0100";
        when x"46f" => qpre <= "0000";
        when x"470" => qpre <= "0000";
        when x"471" => qpre <= "0100";
        when x"472" => qpre <= "0100";
        when x"473" => qpre <= "0000";
        when x"474" => qpre <= "0000";
        when x"475" => qpre <= "0100";
        when x"476" => qpre <= "0100";
        when x"477" => qpre <= "0000";
        when x"478" => qpre <= "0001";
        when x"479" => qpre <= "0101";
        when x"47a" => qpre <= "0101";
        when x"47b" => qpre <= "0001";
        when x"47c" => qpre <= "0000";
        when x"47d" => qpre <= "0000";
        when x"47e" => qpre <= "0000";
        when x"47f" => qpre <= "0000";
        when x"480" => qpre <= "0000";
        when x"481" => qpre <= "0100";
        when x"482" => qpre <= "0100";
        when x"483" => qpre <= "0110";
        when x"484" => qpre <= "0110";
        when x"485" => qpre <= "0110";
        when x"486" => qpre <= "0110";
        when x"487" => qpre <= "0110";
        -- PMICL: disable buck2
        when x"500" => qpre <= "0110";
        when x"501" => qpre <= "0110";
        when x"502" => qpre <= "0110";
        when x"503" => qpre <= "0110";
        when x"504" => qpre <= "0110";
        when x"505" => qpre <= "0100";
        when x"506" => qpre <= "0100";
        when x"507" => qpre <= "0000";
        when x"508" => qpre <= "0010";
        when x"509" => qpre <= "0110";
        when x"50a" => qpre <= "0110";
        when x"50b" => qpre <= "0010";
        when x"50c" => qpre <= "0010";
        when x"50d" => qpre <= "0110";
        when x"50e" => qpre <= "0110";
        when x"50f" => qpre <= "0010";
        when x"510" => qpre <= "0000";
        when x"511" => qpre <= "0100";
        when x"512" => qpre <= "0100";
        when x"513" => qpre <= "0000";
        when x"514" => qpre <= "0000";
        when x"515" => qpre <= "0100";
        when x"516" => qpre <= "0100";
        when x"517" => qpre <= "0000";
        when x"518" => qpre <= "0000";
        when x"519" => qpre <= "0100";
        when x"51a" => qpre <= "0100";
        when x"51b" => qpre <= "0000";
        when x"51c" => qpre <= "0000";
        when x"51d" => qpre <= "0100";
        when x"51e" => qpre <= "0100";
        when x"51f" => qpre <= "0000";
        when x"520" => qpre <= "0000";
        when x"521" => qpre <= "0100";
        when x"522" => qpre <= "0100";
        when x"523" => qpre <= "0000";
        when x"524" => qpre <= "0000";
        when x"525" => qpre <= "0100";
        when x"526" => qpre <= "0100";
        when x"527" => qpre <= "0000";
        when x"528" => qpre <= "0001";
        when x"529" => qpre <= "0101";
        when x"52a" => qpre <= "0101";
        when x"52b" => qpre <= "0001";
        when x"52c" => qpre <= "0000";
        when x"52d" => qpre <= "0000";
        when x"52e" => qpre <= "0000";
        when x"52f" => qpre <= "0000";
        when x"530" => qpre <= "0000";
        when x"531" => qpre <= "0100";
        when x"532" => qpre <= "0100";
        when x"533" => qpre <= "0000";
        when x"534" => qpre <= "0000";
        when x"535" => qpre <= "0100";
        when x"536" => qpre <= "0100";
        when x"537" => qpre <= "0000";
        when x"538" => qpre <= "0000";
        when x"539" => qpre <= "0100";
        when x"53a" => qpre <= "0100";
        when x"53b" => qpre <= "0000";
        when x"53c" => qpre <= "0000";
        when x"53d" => qpre <= "0100";
        when x"53e" => qpre <= "0100";
        when x"53f" => qpre <= "0000";
        when x"540" => qpre <= "0000";
        when x"541" => qpre <= "0100";
        when x"542" => qpre <= "0100";
        when x"543" => qpre <= "0000";
        when x"544" => qpre <= "0010";
        when x"545" => qpre <= "0110";
        when x"546" => qpre <= "0110";
        when x"547" => qpre <= "0010";
        when x"548" => qpre <= "0010";
        when x"549" => qpre <= "0110";
        when x"54a" => qpre <= "0110";
        when x"54b" => qpre <= "0010";
        when x"54c" => qpre <= "0000";
        when x"54d" => qpre <= "0100";
        when x"54e" => qpre <= "0100";
        when x"54f" => qpre <= "0000";
        when x"550" => qpre <= "0001";
        when x"551" => qpre <= "0101";
        when x"552" => qpre <= "0101";
        when x"553" => qpre <= "0001";
        when x"554" => qpre <= "0000";
        when x"555" => qpre <= "0000";
        when x"556" => qpre <= "0000";
        when x"557" => qpre <= "0000";
        when x"558" => qpre <= "0010";
        when x"559" => qpre <= "0110";
        when x"55a" => qpre <= "0110";
        when x"55b" => qpre <= "0010";
        when x"55c" => qpre <= "0010";
        when x"55d" => qpre <= "0110";
        when x"55e" => qpre <= "0110";
        when x"55f" => qpre <= "0010";
        when x"560" => qpre <= "0000";
        when x"561" => qpre <= "0100";
        when x"562" => qpre <= "0100";
        when x"563" => qpre <= "0000";
        when x"564" => qpre <= "0000";
        when x"565" => qpre <= "0100";
        when x"566" => qpre <= "0100";
        when x"567" => qpre <= "0000";
        when x"568" => qpre <= "0010";
        when x"569" => qpre <= "0110";
        when x"56a" => qpre <= "0110";
        when x"56b" => qpre <= "0010";
        when x"56c" => qpre <= "0000";
        when x"56d" => qpre <= "0100";
        when x"56e" => qpre <= "0100";
        when x"56f" => qpre <= "0000";
        when x"570" => qpre <= "0000";
        when x"571" => qpre <= "0100";
        when x"572" => qpre <= "0100";
        when x"573" => qpre <= "0000";
        when x"574" => qpre <= "0000";
        when x"575" => qpre <= "0100";
        when x"576" => qpre <= "0100";
        when x"577" => qpre <= "0000";
        when x"578" => qpre <= "0001";
        when x"579" => qpre <= "0101";
        when x"57a" => qpre <= "0101";
        when x"57b" => qpre <= "0001";
        when x"57c" => qpre <= "0000";
        when x"57d" => qpre <= "0000";
        when x"57e" => qpre <= "0000";
        when x"57f" => qpre <= "0000";
        when x"580" => qpre <= "0000";
        when x"581" => qpre <= "0100";
        when x"582" => qpre <= "0100";
        when x"583" => qpre <= "0110";
        when x"584" => qpre <= "0110";
        when x"585" => qpre <= "0110";
        when x"586" => qpre <= "0110";
        when x"587" => qpre <= "0110";
        -- PMICL: disable buck3
        when x"600" => qpre <= "0110";
        when x"601" => qpre <= "0110";
        when x"602" => qpre <= "0110";
        when x"603" => qpre <= "0110";
        when x"604" => qpre <= "0110";
        when x"605" => qpre <= "0100";
        when x"606" => qpre <= "0100";
        when x"607" => qpre <= "0000";
        when x"608" => qpre <= "0010";
        when x"609" => qpre <= "0110";
        when x"60a" => qpre <= "0110";
        when x"60b" => qpre <= "0010";
        when x"60c" => qpre <= "0010";
        when x"60d" => qpre <= "0110";
        when x"60e" => qpre <= "0110";
        when x"60f" => qpre <= "0010";
        when x"610" => qpre <= "0000";
        when x"611" => qpre <= "0100";
        when x"612" => qpre <= "0100";
        when x"613" => qpre <= "0000";
        when x"614" => qpre <= "0000";
        when x"615" => qpre <= "0100";
        when x"616" => qpre <= "0100";
        when x"617" => qpre <= "0000";
        when x"618" => qpre <= "0000";
        when x"619" => qpre <= "0100";
        when x"61a" => qpre <= "0100";
        when x"61b" => qpre <= "0000";
        when x"61c" => qpre <= "0000";
        when x"61d" => qpre <= "0100";
        when x"61e" => qpre <= "0100";
        when x"61f" => qpre <= "0000";
        when x"620" => qpre <= "0000";
        when x"621" => qpre <= "0100";
        when x"622" => qpre <= "0100";
        when x"623" => qpre <= "0000";
        when x"624" => qpre <= "0000";
        when x"625" => qpre <= "0100";
        when x"626" => qpre <= "0100";
        when x"627" => qpre <= "0000";
        when x"628" => qpre <= "0001";
        when x"629" => qpre <= "0101";
        when x"62a" => qpre <= "0101";
        when x"62b" => qpre <= "0001";
        when x"62c" => qpre <= "0000";
        when x"62d" => qpre <= "0000";
        when x"62e" => qpre <= "0000";
        when x"62f" => qpre <= "0000";
        when x"630" => qpre <= "0000";
        when x"631" => qpre <= "0100";
        when x"632" => qpre <= "0100";
        when x"633" => qpre <= "0000";
        when x"634" => qpre <= "0000";
        when x"635" => qpre <= "0100";
        when x"636" => qpre <= "0100";
        when x"637" => qpre <= "0000";
        when x"638" => qpre <= "0000";
        when x"639" => qpre <= "0100";
        when x"63a" => qpre <= "0100";
        when x"63b" => qpre <= "0000";
        when x"63c" => qpre <= "0000";
        when x"63d" => qpre <= "0100";
        when x"63e" => qpre <= "0100";
        when x"63f" => qpre <= "0000";
        when x"640" => qpre <= "0010";
        when x"641" => qpre <= "0110";
        when x"642" => qpre <= "0110";
        when x"643" => qpre <= "0010";
        when x"644" => qpre <= "0000";
        when x"645" => qpre <= "0100";
        when x"646" => qpre <= "0100";
        when x"647" => qpre <= "0000";
        when x"648" => qpre <= "0000";
        when x"649" => qpre <= "0100";
        when x"64a" => qpre <= "0100";
        when x"64b" => qpre <= "0000";
        when x"64c" => qpre <= "0000";
        when x"64d" => qpre <= "0100";
        when x"64e" => qpre <= "0100";
        when x"64f" => qpre <= "0000";
        when x"650" => qpre <= "0001";
        when x"651" => qpre <= "0101";
        when x"652" => qpre <= "0101";
        when x"653" => qpre <= "0001";
        when x"654" => qpre <= "0000";
        when x"655" => qpre <= "0000";
        when x"656" => qpre <= "0000";
        when x"657" => qpre <= "0000";
        when x"658" => qpre <= "0010";
        when x"659" => qpre <= "0110";
        when x"65a" => qpre <= "0110";
        when x"65b" => qpre <= "0010";
        when x"65c" => qpre <= "0010";
        when x"65d" => qpre <= "0110";
        when x"65e" => qpre <= "0110";
        when x"65f" => qpre <= "0010";
        when x"660" => qpre <= "0000";
        when x"661" => qpre <= "0100";
        when x"662" => qpre <= "0100";
        when x"663" => qpre <= "0000";
        when x"664" => qpre <= "0000";
        when x"665" => qpre <= "0100";
        when x"666" => qpre <= "0100";
        when x"667" => qpre <= "0000";
        when x"668" => qpre <= "0010";
        when x"669" => qpre <= "0110";
        when x"66a" => qpre <= "0110";
        when x"66b" => qpre <= "0010";
        when x"66c" => qpre <= "0000";
        when x"66d" => qpre <= "0100";
        when x"66e" => qpre <= "0100";
        when x"66f" => qpre <= "0000";
        when x"670" => qpre <= "0000";
        when x"671" => qpre <= "0100";
        when x"672" => qpre <= "0100";
        when x"673" => qpre <= "0000";
        when x"674" => qpre <= "0000";
        when x"675" => qpre <= "0100";
        when x"676" => qpre <= "0100";
        when x"677" => qpre <= "0000";
        when x"678" => qpre <= "0001";
        when x"679" => qpre <= "0101";
        when x"67a" => qpre <= "0101";
        when x"67b" => qpre <= "0001";
        when x"67c" => qpre <= "0000";
        when x"67d" => qpre <= "0000";
        when x"67e" => qpre <= "0000";
        when x"67f" => qpre <= "0000";
        when x"680" => qpre <= "0000";
        when x"681" => qpre <= "0100";
        when x"682" => qpre <= "0100";
        when x"683" => qpre <= "0110";
        when x"684" => qpre <= "0110";
        when x"685" => qpre <= "0110";
        when x"686" => qpre <= "0110";
        when x"687" => qpre <= "0110";
        -- PMICL: set buck0 to 1880 mV
        when x"700" => qpre <= "0110";
        when x"701" => qpre <= "0110";
        when x"702" => qpre <= "0110";
        when x"703" => qpre <= "0110";
        when x"704" => qpre <= "0110";
        when x"705" => qpre <= "0100";
        when x"706" => qpre <= "0100";
        when x"707" => qpre <= "0000";
        when x"708" => qpre <= "0010";
        when x"709" => qpre <= "0110";
        when x"70a" => qpre <= "0110";
        when x"70b" => qpre <= "0010";
        when x"70c" => qpre <= "0010";
        when x"70d" => qpre <= "0110";
        when x"70e" => qpre <= "0110";
        when x"70f" => qpre <= "0010";
        when x"710" => qpre <= "0000";
        when x"711" => qpre <= "0100";
        when x"712" => qpre <= "0100";
        when x"713" => qpre <= "0000";
        when x"714" => qpre <= "0000";
        when x"715" => qpre <= "0100";
        when x"716" => qpre <= "0100";
        when x"717" => qpre <= "0000";
        when x"718" => qpre <= "0000";
        when x"719" => qpre <= "0100";
        when x"71a" => qpre <= "0100";
        when x"71b" => qpre <= "0000";
        when x"71c" => qpre <= "0000";
        when x"71d" => qpre <= "0100";
        when x"71e" => qpre <= "0100";
        when x"71f" => qpre <= "0000";
        when x"720" => qpre <= "0000";
        when x"721" => qpre <= "0100";
        when x"722" => qpre <= "0100";
        when x"723" => qpre <= "0000";
        when x"724" => qpre <= "0000";
        when x"725" => qpre <= "0100";
        when x"726" => qpre <= "0100";
        when x"727" => qpre <= "0000";
        when x"728" => qpre <= "0001";
        when x"729" => qpre <= "0101";
        when x"72a" => qpre <= "0101";
        when x"72b" => qpre <= "0001";
        when x"72c" => qpre <= "0000";
        when x"72d" => qpre <= "0000";
        when x"72e" => qpre <= "0000";
        when x"72f" => qpre <= "0000";
        when x"730" => qpre <= "0000";
        when x"731" => qpre <= "0100";
        when x"732" => qpre <= "0100";
        when x"733" => qpre <= "0000";
        when x"734" => qpre <= "0000";
        when x"735" => qpre <= "0100";
        when x"736" => qpre <= "0100";
        when x"737" => qpre <= "0000";
        when x"738" => qpre <= "0000";
        when x"739" => qpre <= "0100";
        when x"73a" => qpre <= "0100";
        when x"73b" => qpre <= "0000";
        when x"73c" => qpre <= "0000";
        when x"73d" => qpre <= "0100";
        when x"73e" => qpre <= "0100";
        when x"73f" => qpre <= "0000";
        when x"740" => qpre <= "0010";
        when x"741" => qpre <= "0110";
        when x"742" => qpre <= "0110";
        when x"743" => qpre <= "0010";
        when x"744" => qpre <= "0000";
        when x"745" => qpre <= "0100";
        when x"746" => qpre <= "0100";
        when x"747" => qpre <= "0000";
        when x"748" => qpre <= "0010";
        when x"749" => qpre <= "0110";
        when x"74a" => qpre <= "0110";
        when x"74b" => qpre <= "0010";
        when x"74c" => qpre <= "0000";
        when x"74d" => qpre <= "0100";
        when x"74e" => qpre <= "0100";
        when x"74f" => qpre <= "0000";
        when x"750" => qpre <= "0001";
        when x"751" => qpre <= "0101";
        when x"752" => qpre <= "0101";
        when x"753" => qpre <= "0001";
        when x"754" => qpre <= "0000";
        when x"755" => qpre <= "0000";
        when x"756" => qpre <= "0000";
        when x"757" => qpre <= "0000";
        when x"758" => qpre <= "0010";
        when x"759" => qpre <= "0110";
        when x"75a" => qpre <= "0110";
        when x"75b" => qpre <= "0010";
        when x"75c" => qpre <= "0000";
        when x"75d" => qpre <= "0100";
        when x"75e" => qpre <= "0100";
        when x"75f" => qpre <= "0000";
        when x"760" => qpre <= "0010";
        when x"761" => qpre <= "0110";
        when x"762" => qpre <= "0110";
        when x"763" => qpre <= "0010";
        when x"764" => qpre <= "0010";
        when x"765" => qpre <= "0110";
        when x"766" => qpre <= "0110";
        when x"767" => qpre <= "0010";
        when x"768" => qpre <= "0000";
        when x"769" => qpre <= "0100";
        when x"76a" => qpre <= "0100";
        when x"76b" => qpre <= "0000";
        when x"76c" => qpre <= "0010";
        when x"76d" => qpre <= "0110";
        when x"76e" => qpre <= "0110";
        when x"76f" => qpre <= "0010";
        when x"770" => qpre <= "0000";
        when x"771" => qpre <= "0100";
        when x"772" => qpre <= "0100";
        when x"773" => qpre <= "0000";
        when x"774" => qpre <= "0010";
        when x"775" => qpre <= "0110";
        when x"776" => qpre <= "0110";
        when x"777" => qpre <= "0010";
        when x"778" => qpre <= "0001";
        when x"779" => qpre <= "0101";
        when x"77a" => qpre <= "0101";
        when x"77b" => qpre <= "0001";
        when x"77c" => qpre <= "0000";
        when x"77d" => qpre <= "0000";
        when x"77e" => qpre <= "0000";
        when x"77f" => qpre <= "0000";
        when x"780" => qpre <= "0000";
        when x"781" => qpre <= "0100";
        when x"782" => qpre <= "0100";
        when x"783" => qpre <= "0110";
        when x"784" => qpre <= "0110";
        when x"785" => qpre <= "0110";
        when x"786" => qpre <= "0110";
        when x"787" => qpre <= "0110";
        -- PMICL: set buck2 to 1480 mV
        when x"800" => qpre <= "0110";
        when x"801" => qpre <= "0110";
        when x"802" => qpre <= "0110";
        when x"803" => qpre <= "0110";
        when x"804" => qpre <= "0110";
        when x"805" => qpre <= "0100";
        when x"806" => qpre <= "0100";
        when x"807" => qpre <= "0000";
        when x"808" => qpre <= "0010";
        when x"809" => qpre <= "0110";
        when x"80a" => qpre <= "0110";
        when x"80b" => qpre <= "0010";
        when x"80c" => qpre <= "0010";
        when x"80d" => qpre <= "0110";
        when x"80e" => qpre <= "0110";
        when x"80f" => qpre <= "0010";
        when x"810" => qpre <= "0000";
        when x"811" => qpre <= "0100";
        when x"812" => qpre <= "0100";
        when x"813" => qpre <= "0000";
        when x"814" => qpre <= "0000";
        when x"815" => qpre <= "0100";
        when x"816" => qpre <= "0100";
        when x"817" => qpre <= "0000";
        when x"818" => qpre <= "0000";
        when x"819" => qpre <= "0100";
        when x"81a" => qpre <= "0100";
        when x"81b" => qpre <= "0000";
        when x"81c" => qpre <= "0000";
        when x"81d" => qpre <= "0100";
        when x"81e" => qpre <= "0100";
        when x"81f" => qpre <= "0000";
        when x"820" => qpre <= "0000";
        when x"821" => qpre <= "0100";
        when x"822" => qpre <= "0100";
        when x"823" => qpre <= "0000";
        when x"824" => qpre <= "0000";
        when x"825" => qpre <= "0100";
        when x"826" => qpre <= "0100";
        when x"827" => qpre <= "0000";
        when x"828" => qpre <= "0001";
        when x"829" => qpre <= "0101";
        when x"82a" => qpre <= "0101";
        when x"82b" => qpre <= "0001";
        when x"82c" => qpre <= "0000";
        when x"82d" => qpre <= "0000";
        when x"82e" => qpre <= "0000";
        when x"82f" => qpre <= "0000";
        when x"830" => qpre <= "0000";
        when x"831" => qpre <= "0100";
        when x"832" => qpre <= "0100";
        when x"833" => qpre <= "0000";
        when x"834" => qpre <= "0000";
        when x"835" => qpre <= "0100";
        when x"836" => qpre <= "0100";
        when x"837" => qpre <= "0000";
        when x"838" => qpre <= "0000";
        when x"839" => qpre <= "0100";
        when x"83a" => qpre <= "0100";
        when x"83b" => qpre <= "0000";
        when x"83c" => qpre <= "0000";
        when x"83d" => qpre <= "0100";
        when x"83e" => qpre <= "0100";
        when x"83f" => qpre <= "0000";
        when x"840" => qpre <= "0010";
        when x"841" => qpre <= "0110";
        when x"842" => qpre <= "0110";
        when x"843" => qpre <= "0010";
        when x"844" => qpre <= "0010";
        when x"845" => qpre <= "0110";
        when x"846" => qpre <= "0110";
        when x"847" => qpre <= "0010";
        when x"848" => qpre <= "0010";
        when x"849" => qpre <= "0110";
        when x"84a" => qpre <= "0110";
        when x"84b" => qpre <= "0010";
        when x"84c" => qpre <= "0000";
        when x"84d" => qpre <= "0100";
        when x"84e" => qpre <= "0100";
        when x"84f" => qpre <= "0000";
        when x"850" => qpre <= "0001";
        when x"851" => qpre <= "0101";
        when x"852" => qpre <= "0101";
        when x"853" => qpre <= "0001";
        when x"854" => qpre <= "0000";
        when x"855" => qpre <= "0000";
        when x"856" => qpre <= "0000";
        when x"857" => qpre <= "0000";
        when x"858" => qpre <= "0010";
        when x"859" => qpre <= "0110";
        when x"85a" => qpre <= "0110";
        when x"85b" => qpre <= "0010";
        when x"85c" => qpre <= "0000";
        when x"85d" => qpre <= "0100";
        when x"85e" => qpre <= "0100";
        when x"85f" => qpre <= "0000";
        when x"860" => qpre <= "0010";
        when x"861" => qpre <= "0110";
        when x"862" => qpre <= "0110";
        when x"863" => qpre <= "0010";
        when x"864" => qpre <= "0000";
        when x"865" => qpre <= "0100";
        when x"866" => qpre <= "0100";
        when x"867" => qpre <= "0000";
        when x"868" => qpre <= "0000";
        when x"869" => qpre <= "0100";
        when x"86a" => qpre <= "0100";
        when x"86b" => qpre <= "0000";
        when x"86c" => qpre <= "0000";
        when x"86d" => qpre <= "0100";
        when x"86e" => qpre <= "0100";
        when x"86f" => qpre <= "0000";
        when x"870" => qpre <= "0000";
        when x"871" => qpre <= "0100";
        when x"872" => qpre <= "0100";
        when x"873" => qpre <= "0000";
        when x"874" => qpre <= "0010";
        when x"875" => qpre <= "0110";
        when x"876" => qpre <= "0110";
        when x"877" => qpre <= "0010";
        when x"878" => qpre <= "0001";
        when x"879" => qpre <= "0101";
        when x"87a" => qpre <= "0101";
        when x"87b" => qpre <= "0001";
        when x"87c" => qpre <= "0000";
        when x"87d" => qpre <= "0000";
        when x"87e" => qpre <= "0000";
        when x"87f" => qpre <= "0000";
        when x"880" => qpre <= "0000";
        when x"881" => qpre <= "0100";
        when x"882" => qpre <= "0100";
        when x"883" => qpre <= "0110";
        when x"884" => qpre <= "0110";
        when x"885" => qpre <= "0110";
        when x"886" => qpre <= "0110";
        when x"887" => qpre <= "0110";
        -- PMICL: set buck3 to 1340 mV
        when x"900" => qpre <= "0110";
        when x"901" => qpre <= "0110";
        when x"902" => qpre <= "0110";
        when x"903" => qpre <= "0110";
        when x"904" => qpre <= "0110";
        when x"905" => qpre <= "0100";
        when x"906" => qpre <= "0100";
        when x"907" => qpre <= "0000";
        when x"908" => qpre <= "0010";
        when x"909" => qpre <= "0110";
        when x"90a" => qpre <= "0110";
        when x"90b" => qpre <= "0010";
        when x"90c" => qpre <= "0010";
        when x"90d" => qpre <= "0110";
        when x"90e" => qpre <= "0110";
        when x"90f" => qpre <= "0010";
        when x"910" => qpre <= "0000";
        when x"911" => qpre <= "0100";
        when x"912" => qpre <= "0100";
        when x"913" => qpre <= "0000";
        when x"914" => qpre <= "0000";
        when x"915" => qpre <= "0100";
        when x"916" => qpre <= "0100";
        when x"917" => qpre <= "0000";
        when x"918" => qpre <= "0000";
        when x"919" => qpre <= "0100";
        when x"91a" => qpre <= "0100";
        when x"91b" => qpre <= "0000";
        when x"91c" => qpre <= "0000";
        when x"91d" => qpre <= "0100";
        when x"91e" => qpre <= "0100";
        when x"91f" => qpre <= "0000";
        when x"920" => qpre <= "0000";
        when x"921" => qpre <= "0100";
        when x"922" => qpre <= "0100";
        when x"923" => qpre <= "0000";
        when x"924" => qpre <= "0000";
        when x"925" => qpre <= "0100";
        when x"926" => qpre <= "0100";
        when x"927" => qpre <= "0000";
        when x"928" => qpre <= "0001";
        when x"929" => qpre <= "0101";
        when x"92a" => qpre <= "0101";
        when x"92b" => qpre <= "0001";
        when x"92c" => qpre <= "0000";
        when x"92d" => qpre <= "0000";
        when x"92e" => qpre <= "0000";
        when x"92f" => qpre <= "0000";
        when x"930" => qpre <= "0000";
        when x"931" => qpre <= "0100";
        when x"932" => qpre <= "0100";
        when x"933" => qpre <= "0000";
        when x"934" => qpre <= "0000";
        when x"935" => qpre <= "0100";
        when x"936" => qpre <= "0100";
        when x"937" => qpre <= "0000";
        when x"938" => qpre <= "0000";
        when x"939" => qpre <= "0100";
        when x"93a" => qpre <= "0100";
        when x"93b" => qpre <= "0000";
        when x"93c" => qpre <= "0010";
        when x"93d" => qpre <= "0110";
        when x"93e" => qpre <= "0110";
        when x"93f" => qpre <= "0010";
        when x"940" => qpre <= "0000";
        when x"941" => qpre <= "0100";
        when x"942" => qpre <= "0100";
        when x"943" => qpre <= "0000";
        when x"944" => qpre <= "0000";
        when x"945" => qpre <= "0100";
        when x"946" => qpre <= "0100";
        when x"947" => qpre <= "0000";
        when x"948" => qpre <= "0000";
        when x"949" => qpre <= "0100";
        when x"94a" => qpre <= "0100";
        when x"94b" => qpre <= "0000";
        when x"94c" => qpre <= "0000";
        when x"94d" => qpre <= "0100";
        when x"94e" => qpre <= "0100";
        when x"94f" => qpre <= "0000";
        when x"950" => qpre <= "0001";
        when x"951" => qpre <= "0101";
        when x"952" => qpre <= "0101";
        when x"953" => qpre <= "0001";
        when x"954" => qpre <= "0000";
        when x"955" => qpre <= "0000";
        when x"956" => qpre <= "0000";
        when x"957" => qpre <= "0000";
        when x"958" => qpre <= "0010";
        when x"959" => qpre <= "0110";
        when x"95a" => qpre <= "0110";
        when x"95b" => qpre <= "0010";
        when x"95c" => qpre <= "0000";
        when x"95d" => qpre <= "0100";
        when x"95e" => qpre <= "0100";
        when x"95f" => qpre <= "0000";
        when x"960" => qpre <= "0000";
        when x"961" => qpre <= "0100";
        when x"962" => qpre <= "0100";
        when x"963" => qpre <= "0000";
        when x"964" => qpre <= "0010";
        when x"965" => qpre <= "0110";
        when x"966" => qpre <= "0110";
        when x"967" => qpre <= "0010";
        when x"968" => qpre <= "0000";
        when x"969" => qpre <= "0100";
        when x"96a" => qpre <= "0100";
        when x"96b" => qpre <= "0000";
        when x"96c" => qpre <= "0000";
        when x"96d" => qpre <= "0100";
        when x"96e" => qpre <= "0100";
        when x"96f" => qpre <= "0000";
        when x"970" => qpre <= "0010";
        when x"971" => qpre <= "0110";
        when x"972" => qpre <= "0110";
        when x"973" => qpre <= "0010";
        when x"974" => qpre <= "0000";
        when x"975" => qpre <= "0100";
        when x"976" => qpre <= "0100";
        when x"977" => qpre <= "0000";
        when x"978" => qpre <= "0001";
        when x"979" => qpre <= "0101";
        when x"97a" => qpre <= "0101";
        when x"97b" => qpre <= "0001";
        when x"97c" => qpre <= "0000";
        when x"97d" => qpre <= "0000";
        when x"97e" => qpre <= "0000";
        when x"97f" => qpre <= "0000";
        when x"980" => qpre <= "0000";
        when x"981" => qpre <= "0100";
        when x"982" => qpre <= "0100";
        when x"983" => qpre <= "0110";
        when x"984" => qpre <= "0110";
        when x"985" => qpre <= "0110";
        when x"986" => qpre <= "0110";
        when x"987" => qpre <= "0110";
        -- delay to make sure PMICF is ready
        -- PMICF: check OTP ID
        when x"b00" => qpre <= "1110";
        when x"b01" => qpre <= "1110";
        when x"b02" => qpre <= "1110";
        when x"b03" => qpre <= "1110";
        when x"b04" => qpre <= "1110";
        when x"b05" => qpre <= "1100";
        when x"b06" => qpre <= "1100";
        when x"b07" => qpre <= "1000";
        when x"b08" => qpre <= "1010";
        when x"b09" => qpre <= "1110";
        when x"b0a" => qpre <= "1110";
        when x"b0b" => qpre <= "1010";
        when x"b0c" => qpre <= "1010";
        when x"b0d" => qpre <= "1110";
        when x"b0e" => qpre <= "1110";
        when x"b0f" => qpre <= "1010";
        when x"b10" => qpre <= "1000";
        when x"b11" => qpre <= "1100";
        when x"b12" => qpre <= "1100";
        when x"b13" => qpre <= "1000";
        when x"b14" => qpre <= "1000";
        when x"b15" => qpre <= "1100";
        when x"b16" => qpre <= "1100";
        when x"b17" => qpre <= "1000";
        when x"b18" => qpre <= "1000";
        when x"b19" => qpre <= "1100";
        when x"b1a" => qpre <= "1100";
        when x"b1b" => qpre <= "1000";
        when x"b1c" => qpre <= "1000";
        when x"b1d" => qpre <= "1100";
        when x"b1e" => qpre <= "1100";
        when x"b1f" => qpre <= "1000";
        when x"b20" => qpre <= "1000";
        when x"b21" => qpre <= "1100";
        when x"b22" => qpre <= "1100";
        when x"b23" => qpre <= "1000";
        when x"b24" => qpre <= "1000";
        when x"b25" => qpre <= "1100";
        when x"b26" => qpre <= "1100";
        when x"b27" => qpre <= "1000";
        when x"b28" => qpre <= "1001";
        when x"b29" => qpre <= "1101";
        when x"b2a" => qpre <= "1101";
        when x"b2b" => qpre <= "1001";
        when x"b2c" => qpre <= "1000";
        when x"b2d" => qpre <= "1000";
        when x"b2e" => qpre <= "1000";
        when x"b2f" => qpre <= "1000";
        when x"b30" => qpre <= "1000";
        when x"b31" => qpre <= "1100";
        when x"b32" => qpre <= "1100";
        when x"b33" => qpre <= "1000";
        when x"b34" => qpre <= "1000";
        when x"b35" => qpre <= "1100";
        when x"b36" => qpre <= "1100";
        when x"b37" => qpre <= "1000";
        when x"b38" => qpre <= "1000";
        when x"b39" => qpre <= "1100";
        when x"b3a" => qpre <= "1100";
        when x"b3b" => qpre <= "1000";
        when x"b3c" => qpre <= "1000";
        when x"b3d" => qpre <= "1100";
        when x"b3e" => qpre <= "1100";
        when x"b3f" => qpre <= "1000";
        when x"b40" => qpre <= "1000";
        when x"b41" => qpre <= "1100";
        when x"b42" => qpre <= "1100";
        when x"b43" => qpre <= "1000";
        when x"b44" => qpre <= "1000";
        when x"b45" => qpre <= "1100";
        when x"b46" => qpre <= "1100";
        when x"b47" => qpre <= "1000";
        when x"b48" => qpre <= "1000";
        when x"b49" => qpre <= "1100";
        when x"b4a" => qpre <= "1100";
        when x"b4b" => qpre <= "1000";
        when x"b4c" => qpre <= "1010";
        when x"b4d" => qpre <= "1110";
        when x"b4e" => qpre <= "1110";
        when x"b4f" => qpre <= "1010";
        when x"b50" => qpre <= "1001";
        when x"b51" => qpre <= "1101";
        when x"b52" => qpre <= "1101";
        when x"b53" => qpre <= "1001";
        when x"b54" => qpre <= "1010";
        when x"b55" => qpre <= "1110";
        when x"b56" => qpre <= "1100";
        when x"b57" => qpre <= "1000";
        when x"b58" => qpre <= "1010";
        when x"b59" => qpre <= "1110";
        when x"b5a" => qpre <= "1110";
        when x"b5b" => qpre <= "1010";
        when x"b5c" => qpre <= "1010";
        when x"b5d" => qpre <= "1110";
        when x"b5e" => qpre <= "1110";
        when x"b5f" => qpre <= "1010";
        when x"b60" => qpre <= "1000";
        when x"b61" => qpre <= "1100";
        when x"b62" => qpre <= "1100";
        when x"b63" => qpre <= "1000";
        when x"b64" => qpre <= "1000";
        when x"b65" => qpre <= "1100";
        when x"b66" => qpre <= "1100";
        when x"b67" => qpre <= "1000";
        when x"b68" => qpre <= "1000";
        when x"b69" => qpre <= "1100";
        when x"b6a" => qpre <= "1100";
        when x"b6b" => qpre <= "1000";
        when x"b6c" => qpre <= "1000";
        when x"b6d" => qpre <= "1100";
        when x"b6e" => qpre <= "1100";
        when x"b6f" => qpre <= "1000";
        when x"b70" => qpre <= "1000";
        when x"b71" => qpre <= "1100";
        when x"b72" => qpre <= "1100";
        when x"b73" => qpre <= "1000";
        when x"b74" => qpre <= "1010";
        when x"b75" => qpre <= "1110";
        when x"b76" => qpre <= "1110";
        when x"b77" => qpre <= "1010";
        when x"b78" => qpre <= "1001";
        when x"b79" => qpre <= "1101";
        when x"b7a" => qpre <= "1101";
        when x"b7b" => qpre <= "1001";
        when x"b7c" => qpre <= "1000";
        when x"b7d" => qpre <= "1000";
        when x"b7e" => qpre <= "1000";
        when x"b7f" => qpre <= "1000";
        when x"b80" => qpre <= "1011";
        when x"b81" => qpre <= "1111";
        when x"b82" => qpre <= "1111";
        when x"b83" => qpre <= "1011";
        when x"b84" => qpre <= "1011";
        when x"b85" => qpre <= "1111";
        when x"b86" => qpre <= "1111";
        when x"b87" => qpre <= "1011";
        when x"b88" => qpre <= "1011";
        when x"b89" => qpre <= "1111";
        when x"b8a" => qpre <= "1111";
        when x"b8b" => qpre <= "1011";
        when x"b8c" => qpre <= "1001";
        when x"b8d" => qpre <= "1101";
        when x"b8e" => qpre <= "1101";
        when x"b8f" => qpre <= "1001";
        when x"b90" => qpre <= "1001";
        when x"b91" => qpre <= "1101";
        when x"b92" => qpre <= "1101";
        when x"b93" => qpre <= "1001";
        when x"b94" => qpre <= "1001";
        when x"b95" => qpre <= "1101";
        when x"b96" => qpre <= "1101";
        when x"b97" => qpre <= "1001";
        when x"b98" => qpre <= "1001";
        when x"b99" => qpre <= "1101";
        when x"b9a" => qpre <= "1101";
        when x"b9b" => qpre <= "1001";
        when x"b9c" => qpre <= "1001";
        when x"b9d" => qpre <= "1101";
        when x"b9e" => qpre <= "1101";
        when x"b9f" => qpre <= "1001";
        when x"ba0" => qpre <= "1010";
        when x"ba1" => qpre <= "1110";
        when x"ba2" => qpre <= "1110";
        when x"ba3" => qpre <= "1010";
        when x"ba4" => qpre <= "1000";
        when x"ba5" => qpre <= "1000";
        when x"ba6" => qpre <= "1000";
        when x"ba7" => qpre <= "1000";
        when x"ba8" => qpre <= "1000";
        when x"ba9" => qpre <= "1100";
        when x"baa" => qpre <= "1100";
        when x"bab" => qpre <= "1110";
        when x"bac" => qpre <= "1110";
        when x"bad" => qpre <= "1110";
        when x"bae" => qpre <= "1110";
        when x"baf" => qpre <= "1110";
        -- PMICL: enable buck0
        when x"c00" => qpre <= "0110";
        when x"c01" => qpre <= "0110";
        when x"c02" => qpre <= "0110";
        when x"c03" => qpre <= "0110";
        when x"c04" => qpre <= "0110";
        when x"c05" => qpre <= "0100";
        when x"c06" => qpre <= "0100";
        when x"c07" => qpre <= "0000";
        when x"c08" => qpre <= "0010";
        when x"c09" => qpre <= "0110";
        when x"c0a" => qpre <= "0110";
        when x"c0b" => qpre <= "0010";
        when x"c0c" => qpre <= "0010";
        when x"c0d" => qpre <= "0110";
        when x"c0e" => qpre <= "0110";
        when x"c0f" => qpre <= "0010";
        when x"c10" => qpre <= "0000";
        when x"c11" => qpre <= "0100";
        when x"c12" => qpre <= "0100";
        when x"c13" => qpre <= "0000";
        when x"c14" => qpre <= "0000";
        when x"c15" => qpre <= "0100";
        when x"c16" => qpre <= "0100";
        when x"c17" => qpre <= "0000";
        when x"c18" => qpre <= "0000";
        when x"c19" => qpre <= "0100";
        when x"c1a" => qpre <= "0100";
        when x"c1b" => qpre <= "0000";
        when x"c1c" => qpre <= "0000";
        when x"c1d" => qpre <= "0100";
        when x"c1e" => qpre <= "0100";
        when x"c1f" => qpre <= "0000";
        when x"c20" => qpre <= "0000";
        when x"c21" => qpre <= "0100";
        when x"c22" => qpre <= "0100";
        when x"c23" => qpre <= "0000";
        when x"c24" => qpre <= "0000";
        when x"c25" => qpre <= "0100";
        when x"c26" => qpre <= "0100";
        when x"c27" => qpre <= "0000";
        when x"c28" => qpre <= "0001";
        when x"c29" => qpre <= "0101";
        when x"c2a" => qpre <= "0101";
        when x"c2b" => qpre <= "0001";
        when x"c2c" => qpre <= "0000";
        when x"c2d" => qpre <= "0000";
        when x"c2e" => qpre <= "0000";
        when x"c2f" => qpre <= "0000";
        when x"c30" => qpre <= "0000";
        when x"c31" => qpre <= "0100";
        when x"c32" => qpre <= "0100";
        when x"c33" => qpre <= "0000";
        when x"c34" => qpre <= "0000";
        when x"c35" => qpre <= "0100";
        when x"c36" => qpre <= "0100";
        when x"c37" => qpre <= "0000";
        when x"c38" => qpre <= "0000";
        when x"c39" => qpre <= "0100";
        when x"c3a" => qpre <= "0100";
        when x"c3b" => qpre <= "0000";
        when x"c3c" => qpre <= "0000";
        when x"c3d" => qpre <= "0100";
        when x"c3e" => qpre <= "0100";
        when x"c3f" => qpre <= "0000";
        when x"c40" => qpre <= "0000";
        when x"c41" => qpre <= "0100";
        when x"c42" => qpre <= "0100";
        when x"c43" => qpre <= "0000";
        when x"c44" => qpre <= "0000";
        when x"c45" => qpre <= "0100";
        when x"c46" => qpre <= "0100";
        when x"c47" => qpre <= "0000";
        when x"c48" => qpre <= "0010";
        when x"c49" => qpre <= "0110";
        when x"c4a" => qpre <= "0110";
        when x"c4b" => qpre <= "0010";
        when x"c4c" => qpre <= "0000";
        when x"c4d" => qpre <= "0100";
        when x"c4e" => qpre <= "0100";
        when x"c4f" => qpre <= "0000";
        when x"c50" => qpre <= "0001";
        when x"c51" => qpre <= "0101";
        when x"c52" => qpre <= "0101";
        when x"c53" => qpre <= "0001";
        when x"c54" => qpre <= "0000";
        when x"c55" => qpre <= "0000";
        when x"c56" => qpre <= "0000";
        when x"c57" => qpre <= "0000";
        when x"c58" => qpre <= "0010";
        when x"c59" => qpre <= "0110";
        when x"c5a" => qpre <= "0110";
        when x"c5b" => qpre <= "0010";
        when x"c5c" => qpre <= "0000";
        when x"c5d" => qpre <= "0100";
        when x"c5e" => qpre <= "0100";
        when x"c5f" => qpre <= "0000";
        when x"c60" => qpre <= "0000";
        when x"c61" => qpre <= "0100";
        when x"c62" => qpre <= "0100";
        when x"c63" => qpre <= "0000";
        when x"c64" => qpre <= "0000";
        when x"c65" => qpre <= "0100";
        when x"c66" => qpre <= "0100";
        when x"c67" => qpre <= "0000";
        when x"c68" => qpre <= "0010";
        when x"c69" => qpre <= "0110";
        when x"c6a" => qpre <= "0110";
        when x"c6b" => qpre <= "0010";
        when x"c6c" => qpre <= "0000";
        when x"c6d" => qpre <= "0100";
        when x"c6e" => qpre <= "0100";
        when x"c6f" => qpre <= "0000";
        when x"c70" => qpre <= "0000";
        when x"c71" => qpre <= "0100";
        when x"c72" => qpre <= "0100";
        when x"c73" => qpre <= "0000";
        when x"c74" => qpre <= "0000";
        when x"c75" => qpre <= "0100";
        when x"c76" => qpre <= "0100";
        when x"c77" => qpre <= "0000";
        when x"c78" => qpre <= "0001";
        when x"c79" => qpre <= "0101";
        when x"c7a" => qpre <= "0101";
        when x"c7b" => qpre <= "0001";
        when x"c7c" => qpre <= "0000";
        when x"c7d" => qpre <= "0000";
        when x"c7e" => qpre <= "0000";
        when x"c7f" => qpre <= "0000";
        when x"c80" => qpre <= "0000";
        when x"c81" => qpre <= "0100";
        when x"c82" => qpre <= "0100";
        when x"c83" => qpre <= "0110";
        when x"c84" => qpre <= "0110";
        when x"c85" => qpre <= "0110";
        when x"c86" => qpre <= "0110";
        when x"c87" => qpre <= "0110";
        -- PMICL: enable buck2
        when x"d00" => qpre <= "0110";
        when x"d01" => qpre <= "0110";
        when x"d02" => qpre <= "0110";
        when x"d03" => qpre <= "0110";
        when x"d04" => qpre <= "0110";
        when x"d05" => qpre <= "0100";
        when x"d06" => qpre <= "0100";
        when x"d07" => qpre <= "0000";
        when x"d08" => qpre <= "0010";
        when x"d09" => qpre <= "0110";
        when x"d0a" => qpre <= "0110";
        when x"d0b" => qpre <= "0010";
        when x"d0c" => qpre <= "0010";
        when x"d0d" => qpre <= "0110";
        when x"d0e" => qpre <= "0110";
        when x"d0f" => qpre <= "0010";
        when x"d10" => qpre <= "0000";
        when x"d11" => qpre <= "0100";
        when x"d12" => qpre <= "0100";
        when x"d13" => qpre <= "0000";
        when x"d14" => qpre <= "0000";
        when x"d15" => qpre <= "0100";
        when x"d16" => qpre <= "0100";
        when x"d17" => qpre <= "0000";
        when x"d18" => qpre <= "0000";
        when x"d19" => qpre <= "0100";
        when x"d1a" => qpre <= "0100";
        when x"d1b" => qpre <= "0000";
        when x"d1c" => qpre <= "0000";
        when x"d1d" => qpre <= "0100";
        when x"d1e" => qpre <= "0100";
        when x"d1f" => qpre <= "0000";
        when x"d20" => qpre <= "0000";
        when x"d21" => qpre <= "0100";
        when x"d22" => qpre <= "0100";
        when x"d23" => qpre <= "0000";
        when x"d24" => qpre <= "0000";
        when x"d25" => qpre <= "0100";
        when x"d26" => qpre <= "0100";
        when x"d27" => qpre <= "0000";
        when x"d28" => qpre <= "0001";
        when x"d29" => qpre <= "0101";
        when x"d2a" => qpre <= "0101";
        when x"d2b" => qpre <= "0001";
        when x"d2c" => qpre <= "0000";
        when x"d2d" => qpre <= "0000";
        when x"d2e" => qpre <= "0000";
        when x"d2f" => qpre <= "0000";
        when x"d30" => qpre <= "0000";
        when x"d31" => qpre <= "0100";
        when x"d32" => qpre <= "0100";
        when x"d33" => qpre <= "0000";
        when x"d34" => qpre <= "0000";
        when x"d35" => qpre <= "0100";
        when x"d36" => qpre <= "0100";
        when x"d37" => qpre <= "0000";
        when x"d38" => qpre <= "0000";
        when x"d39" => qpre <= "0100";
        when x"d3a" => qpre <= "0100";
        when x"d3b" => qpre <= "0000";
        when x"d3c" => qpre <= "0000";
        when x"d3d" => qpre <= "0100";
        when x"d3e" => qpre <= "0100";
        when x"d3f" => qpre <= "0000";
        when x"d40" => qpre <= "0000";
        when x"d41" => qpre <= "0100";
        when x"d42" => qpre <= "0100";
        when x"d43" => qpre <= "0000";
        when x"d44" => qpre <= "0010";
        when x"d45" => qpre <= "0110";
        when x"d46" => qpre <= "0110";
        when x"d47" => qpre <= "0010";
        when x"d48" => qpre <= "0010";
        when x"d49" => qpre <= "0110";
        when x"d4a" => qpre <= "0110";
        when x"d4b" => qpre <= "0010";
        when x"d4c" => qpre <= "0000";
        when x"d4d" => qpre <= "0100";
        when x"d4e" => qpre <= "0100";
        when x"d4f" => qpre <= "0000";
        when x"d50" => qpre <= "0001";
        when x"d51" => qpre <= "0101";
        when x"d52" => qpre <= "0101";
        when x"d53" => qpre <= "0001";
        when x"d54" => qpre <= "0000";
        when x"d55" => qpre <= "0000";
        when x"d56" => qpre <= "0000";
        when x"d57" => qpre <= "0000";
        when x"d58" => qpre <= "0010";
        when x"d59" => qpre <= "0110";
        when x"d5a" => qpre <= "0110";
        when x"d5b" => qpre <= "0010";
        when x"d5c" => qpre <= "0000";
        when x"d5d" => qpre <= "0100";
        when x"d5e" => qpre <= "0100";
        when x"d5f" => qpre <= "0000";
        when x"d60" => qpre <= "0000";
        when x"d61" => qpre <= "0100";
        when x"d62" => qpre <= "0100";
        when x"d63" => qpre <= "0000";
        when x"d64" => qpre <= "0000";
        when x"d65" => qpre <= "0100";
        when x"d66" => qpre <= "0100";
        when x"d67" => qpre <= "0000";
        when x"d68" => qpre <= "0010";
        when x"d69" => qpre <= "0110";
        when x"d6a" => qpre <= "0110";
        when x"d6b" => qpre <= "0010";
        when x"d6c" => qpre <= "0000";
        when x"d6d" => qpre <= "0100";
        when x"d6e" => qpre <= "0100";
        when x"d6f" => qpre <= "0000";
        when x"d70" => qpre <= "0000";
        when x"d71" => qpre <= "0100";
        when x"d72" => qpre <= "0100";
        when x"d73" => qpre <= "0000";
        when x"d74" => qpre <= "0000";
        when x"d75" => qpre <= "0100";
        when x"d76" => qpre <= "0100";
        when x"d77" => qpre <= "0000";
        when x"d78" => qpre <= "0001";
        when x"d79" => qpre <= "0101";
        when x"d7a" => qpre <= "0101";
        when x"d7b" => qpre <= "0001";
        when x"d7c" => qpre <= "0000";
        when x"d7d" => qpre <= "0000";
        when x"d7e" => qpre <= "0000";
        when x"d7f" => qpre <= "0000";
        when x"d80" => qpre <= "0000";
        when x"d81" => qpre <= "0100";
        when x"d82" => qpre <= "0100";
        when x"d83" => qpre <= "0110";
        when x"d84" => qpre <= "0110";
        when x"d85" => qpre <= "0110";
        when x"d86" => qpre <= "0110";
        when x"d87" => qpre <= "0110";
        -- PMICL: enable buck3
        when x"e00" => qpre <= "0110";
        when x"e01" => qpre <= "0110";
        when x"e02" => qpre <= "0110";
        when x"e03" => qpre <= "0110";
        when x"e04" => qpre <= "0110";
        when x"e05" => qpre <= "0100";
        when x"e06" => qpre <= "0100";
        when x"e07" => qpre <= "0000";
        when x"e08" => qpre <= "0010";
        when x"e09" => qpre <= "0110";
        when x"e0a" => qpre <= "0110";
        when x"e0b" => qpre <= "0010";
        when x"e0c" => qpre <= "0010";
        when x"e0d" => qpre <= "0110";
        when x"e0e" => qpre <= "0110";
        when x"e0f" => qpre <= "0010";
        when x"e10" => qpre <= "0000";
        when x"e11" => qpre <= "0100";
        when x"e12" => qpre <= "0100";
        when x"e13" => qpre <= "0000";
        when x"e14" => qpre <= "0000";
        when x"e15" => qpre <= "0100";
        when x"e16" => qpre <= "0100";
        when x"e17" => qpre <= "0000";
        when x"e18" => qpre <= "0000";
        when x"e19" => qpre <= "0100";
        when x"e1a" => qpre <= "0100";
        when x"e1b" => qpre <= "0000";
        when x"e1c" => qpre <= "0000";
        when x"e1d" => qpre <= "0100";
        when x"e1e" => qpre <= "0100";
        when x"e1f" => qpre <= "0000";
        when x"e20" => qpre <= "0000";
        when x"e21" => qpre <= "0100";
        when x"e22" => qpre <= "0100";
        when x"e23" => qpre <= "0000";
        when x"e24" => qpre <= "0000";
        when x"e25" => qpre <= "0100";
        when x"e26" => qpre <= "0100";
        when x"e27" => qpre <= "0000";
        when x"e28" => qpre <= "0001";
        when x"e29" => qpre <= "0101";
        when x"e2a" => qpre <= "0101";
        when x"e2b" => qpre <= "0001";
        when x"e2c" => qpre <= "0000";
        when x"e2d" => qpre <= "0000";
        when x"e2e" => qpre <= "0000";
        when x"e2f" => qpre <= "0000";
        when x"e30" => qpre <= "0000";
        when x"e31" => qpre <= "0100";
        when x"e32" => qpre <= "0100";
        when x"e33" => qpre <= "0000";
        when x"e34" => qpre <= "0000";
        when x"e35" => qpre <= "0100";
        when x"e36" => qpre <= "0100";
        when x"e37" => qpre <= "0000";
        when x"e38" => qpre <= "0000";
        when x"e39" => qpre <= "0100";
        when x"e3a" => qpre <= "0100";
        when x"e3b" => qpre <= "0000";
        when x"e3c" => qpre <= "0000";
        when x"e3d" => qpre <= "0100";
        when x"e3e" => qpre <= "0100";
        when x"e3f" => qpre <= "0000";
        when x"e40" => qpre <= "0010";
        when x"e41" => qpre <= "0110";
        when x"e42" => qpre <= "0110";
        when x"e43" => qpre <= "0010";
        when x"e44" => qpre <= "0000";
        when x"e45" => qpre <= "0100";
        when x"e46" => qpre <= "0100";
        when x"e47" => qpre <= "0000";
        when x"e48" => qpre <= "0000";
        when x"e49" => qpre <= "0100";
        when x"e4a" => qpre <= "0100";
        when x"e4b" => qpre <= "0000";
        when x"e4c" => qpre <= "0000";
        when x"e4d" => qpre <= "0100";
        when x"e4e" => qpre <= "0100";
        when x"e4f" => qpre <= "0000";
        when x"e50" => qpre <= "0001";
        when x"e51" => qpre <= "0101";
        when x"e52" => qpre <= "0101";
        when x"e53" => qpre <= "0001";
        when x"e54" => qpre <= "0000";
        when x"e55" => qpre <= "0000";
        when x"e56" => qpre <= "0000";
        when x"e57" => qpre <= "0000";
        when x"e58" => qpre <= "0010";
        when x"e59" => qpre <= "0110";
        when x"e5a" => qpre <= "0110";
        when x"e5b" => qpre <= "0010";
        when x"e5c" => qpre <= "0000";
        when x"e5d" => qpre <= "0100";
        when x"e5e" => qpre <= "0100";
        when x"e5f" => qpre <= "0000";
        when x"e60" => qpre <= "0000";
        when x"e61" => qpre <= "0100";
        when x"e62" => qpre <= "0100";
        when x"e63" => qpre <= "0000";
        when x"e64" => qpre <= "0000";
        when x"e65" => qpre <= "0100";
        when x"e66" => qpre <= "0100";
        when x"e67" => qpre <= "0000";
        when x"e68" => qpre <= "0010";
        when x"e69" => qpre <= "0110";
        when x"e6a" => qpre <= "0110";
        when x"e6b" => qpre <= "0010";
        when x"e6c" => qpre <= "0000";
        when x"e6d" => qpre <= "0100";
        when x"e6e" => qpre <= "0100";
        when x"e6f" => qpre <= "0000";
        when x"e70" => qpre <= "0000";
        when x"e71" => qpre <= "0100";
        when x"e72" => qpre <= "0100";
        when x"e73" => qpre <= "0000";
        when x"e74" => qpre <= "0000";
        when x"e75" => qpre <= "0100";
        when x"e76" => qpre <= "0100";
        when x"e77" => qpre <= "0000";
        when x"e78" => qpre <= "0001";
        when x"e79" => qpre <= "0101";
        when x"e7a" => qpre <= "0101";
        when x"e7b" => qpre <= "0001";
        when x"e7c" => qpre <= "0000";
        when x"e7d" => qpre <= "0000";
        when x"e7e" => qpre <= "0000";
        when x"e7f" => qpre <= "0000";
        when x"e80" => qpre <= "0000";
        when x"e81" => qpre <= "0100";
        when x"e82" => qpre <= "0100";
        when x"e83" => qpre <= "0110";
        when x"e84" => qpre <= "0110";
        when x"e85" => qpre <= "0110";
        when x"e86" => qpre <= "0110";
        when x"e87" => qpre <= "0110";
        -- PMICF: set buck1 to 1800 mV
        when x"f00" => qpre <= "1110";
        when x"f01" => qpre <= "1110";
        when x"f02" => qpre <= "1110";
        when x"f03" => qpre <= "1110";
        when x"f04" => qpre <= "1110";
        when x"f05" => qpre <= "1100";
        when x"f06" => qpre <= "1100";
        when x"f07" => qpre <= "1000";
        when x"f08" => qpre <= "1010";
        when x"f09" => qpre <= "1110";
        when x"f0a" => qpre <= "1110";
        when x"f0b" => qpre <= "1010";
        when x"f0c" => qpre <= "1010";
        when x"f0d" => qpre <= "1110";
        when x"f0e" => qpre <= "1110";
        when x"f0f" => qpre <= "1010";
        when x"f10" => qpre <= "1000";
        when x"f11" => qpre <= "1100";
        when x"f12" => qpre <= "1100";
        when x"f13" => qpre <= "1000";
        when x"f14" => qpre <= "1000";
        when x"f15" => qpre <= "1100";
        when x"f16" => qpre <= "1100";
        when x"f17" => qpre <= "1000";
        when x"f18" => qpre <= "1000";
        when x"f19" => qpre <= "1100";
        when x"f1a" => qpre <= "1100";
        when x"f1b" => qpre <= "1000";
        when x"f1c" => qpre <= "1000";
        when x"f1d" => qpre <= "1100";
        when x"f1e" => qpre <= "1100";
        when x"f1f" => qpre <= "1000";
        when x"f20" => qpre <= "1000";
        when x"f21" => qpre <= "1100";
        when x"f22" => qpre <= "1100";
        when x"f23" => qpre <= "1000";
        when x"f24" => qpre <= "1000";
        when x"f25" => qpre <= "1100";
        when x"f26" => qpre <= "1100";
        when x"f27" => qpre <= "1000";
        when x"f28" => qpre <= "1001";
        when x"f29" => qpre <= "1101";
        when x"f2a" => qpre <= "1101";
        when x"f2b" => qpre <= "1001";
        when x"f2c" => qpre <= "1000";
        when x"f2d" => qpre <= "1000";
        when x"f2e" => qpre <= "1000";
        when x"f2f" => qpre <= "1000";
        when x"f30" => qpre <= "1000";
        when x"f31" => qpre <= "1100";
        when x"f32" => qpre <= "1100";
        when x"f33" => qpre <= "1000";
        when x"f34" => qpre <= "1000";
        when x"f35" => qpre <= "1100";
        when x"f36" => qpre <= "1100";
        when x"f37" => qpre <= "1000";
        when x"f38" => qpre <= "1000";
        when x"f39" => qpre <= "1100";
        when x"f3a" => qpre <= "1100";
        when x"f3b" => qpre <= "1000";
        when x"f3c" => qpre <= "1000";
        when x"f3d" => qpre <= "1100";
        when x"f3e" => qpre <= "1100";
        when x"f3f" => qpre <= "1000";
        when x"f40" => qpre <= "1010";
        when x"f41" => qpre <= "1110";
        when x"f42" => qpre <= "1110";
        when x"f43" => qpre <= "1010";
        when x"f44" => qpre <= "1010";
        when x"f45" => qpre <= "1110";
        when x"f46" => qpre <= "1110";
        when x"f47" => qpre <= "1010";
        when x"f48" => qpre <= "1000";
        when x"f49" => qpre <= "1100";
        when x"f4a" => qpre <= "1100";
        when x"f4b" => qpre <= "1000";
        when x"f4c" => qpre <= "1000";
        when x"f4d" => qpre <= "1100";
        when x"f4e" => qpre <= "1100";
        when x"f4f" => qpre <= "1000";
        when x"f50" => qpre <= "1001";
        when x"f51" => qpre <= "1101";
        when x"f52" => qpre <= "1101";
        when x"f53" => qpre <= "1001";
        when x"f54" => qpre <= "1000";
        when x"f55" => qpre <= "1000";
        when x"f56" => qpre <= "1000";
        when x"f57" => qpre <= "1000";
        when x"f58" => qpre <= "1010";
        when x"f59" => qpre <= "1110";
        when x"f5a" => qpre <= "1110";
        when x"f5b" => qpre <= "1010";
        when x"f5c" => qpre <= "1000";
        when x"f5d" => qpre <= "1100";
        when x"f5e" => qpre <= "1100";
        when x"f5f" => qpre <= "1000";
        when x"f60" => qpre <= "1010";
        when x"f61" => qpre <= "1110";
        when x"f62" => qpre <= "1110";
        when x"f63" => qpre <= "1010";
        when x"f64" => qpre <= "1010";
        when x"f65" => qpre <= "1110";
        when x"f66" => qpre <= "1110";
        when x"f67" => qpre <= "1010";
        when x"f68" => qpre <= "1000";
        when x"f69" => qpre <= "1100";
        when x"f6a" => qpre <= "1100";
        when x"f6b" => qpre <= "1000";
        when x"f6c" => qpre <= "1000";
        when x"f6d" => qpre <= "1100";
        when x"f6e" => qpre <= "1100";
        when x"f6f" => qpre <= "1000";
        when x"f70" => qpre <= "1000";
        when x"f71" => qpre <= "1100";
        when x"f72" => qpre <= "1100";
        when x"f73" => qpre <= "1000";
        when x"f74" => qpre <= "1010";
        when x"f75" => qpre <= "1110";
        when x"f76" => qpre <= "1110";
        when x"f77" => qpre <= "1010";
        when x"f78" => qpre <= "1001";
        when x"f79" => qpre <= "1101";
        when x"f7a" => qpre <= "1101";
        when x"f7b" => qpre <= "1001";
        when x"f7c" => qpre <= "1000";
        when x"f7d" => qpre <= "1000";
        when x"f7e" => qpre <= "1000";
        when x"f7f" => qpre <= "1000";
        when x"f80" => qpre <= "1000";
        when x"f81" => qpre <= "1100";
        when x"f82" => qpre <= "1100";
        when x"f83" => qpre <= "1110";
        when x"f84" => qpre <= "1110";
        when x"f85" => qpre <= "1110";
        when x"f86" => qpre <= "1110";
        when x"f87" => qpre <= "1110";
        -- idle and final state
        when others => qpre <= "1110";
      end case;

      Q <= qpre;

    end if;
  end process;

end architecture imp;


